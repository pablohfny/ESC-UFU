/* testbench para DMux8Way16 */
/* ordem de portas: a, b, c, d, e, f, g, h, in, sel */
/* input [15:0] in; input [2:0] sel; */
/* output [15:0] a; output [15:0] b; output [15:0] c; output [15:0] d; output [15:0] e; output [15:0] f; output [15:0] g; output [15:0] h; */

`include "DMux8Way16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_DMux8Way16;
    reg [15:0] in;
    reg [2:0] sel;
    wire [15:0] a;
    wire [15:0] b;
    wire [15:0] c;
    wire [15:0] d;
    wire [15:0] e;
    wire [15:0] f;
    wire [15:0] g;
    wire [15:0] h;

    DMux8Way16 mymodule(a, b, c, d, e, f, g, h, in, sel);
    
    initial
    begin
        $dumpfile("tb_DMux8Way16.vcd");
        $dumpvars(0, tb_DMux8Way16);

        in = 16'b0000000000000000; sel = 3'b000; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0000010101000110; sel = 3'b000; #1;
         `assert(a, 16'b0000010101000110) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0000011001011000; sel = 3'b110; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000011001011000) `assert(h, 16'b0000000000000000)
        in = 16'b0000111111111100; sel = 3'b101; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000111111111100) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0001000010111110; sel = 3'b110; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0001000010111110) `assert(h, 16'b0000000000000000)
        in = 16'b0001001101100001; sel = 3'b000; #1;
         `assert(a, 16'b0001001101100001) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0001011101101010; sel = 3'b000; #1;
         `assert(a, 16'b0001011101101010) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0001100011011100; sel = 3'b101; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0001100011011100) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0010000111011111; sel = 3'b100; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0010000111011111) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0011000101110111; sel = 3'b011; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0011000101110111) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0100001010001101; sel = 3'b001; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0100001010001101) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0100110011110010; sel = 3'b111; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0100110011110010)
        in = 16'b0101011000001010; sel = 3'b101; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0101011000001010) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0101100001111001; sel = 3'b001; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0101100001111001) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b0110000000111110; sel = 3'b111; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0110000000111110)
        in = 16'b0111100110000100; sel = 3'b110; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0111100110000100) `assert(h, 16'b0000000000000000)
        in = 16'b0111111110110001; sel = 3'b010; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0111111110110001) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1000010111000010; sel = 3'b010; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b1000010111000010) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1000011010111100; sel = 3'b010; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b1000011010111100) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1000111101101000; sel = 3'b101; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b1000111101101000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1001100001100001; sel = 3'b000; #1;
         `assert(a, 16'b1001100001100001) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1001110110111010; sel = 3'b011; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1001110110111010) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1011101110011100; sel = 3'b011; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1011101110011100) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1100010011110100; sel = 3'b101; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b1100010011110100) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1100101001010000; sel = 3'b010; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b1100101001010000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1101100101101000; sel = 3'b110; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b1101100101101000) `assert(h, 16'b0000000000000000)
        in = 16'b1110100100011001; sel = 3'b100; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b1110100100011001) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1111010010111010; sel = 3'b110; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b1111010010111010) `assert(h, 16'b0000000000000000)
        in = 16'b1111100100001100; sel = 3'b101; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b1111100100001100) `assert(g, 16'b0000000000000000) `assert(h, 16'b0000000000000000)
        in = 16'b1111111111111111; sel = 3'b111; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000) `assert(e, 16'b0000000000000000) `assert(f, 16'b0000000000000000) `assert(g, 16'b0000000000000000) `assert(h, 16'b1111111111111111)

    end
endmodule