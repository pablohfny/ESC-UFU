/* testbench para Or16 */
/* ordem de portas: out, a, b */
/* input [15:0] a; input [15:0] b; */
/* output [15:0] out; */

`include "Or16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_Or16;
    reg [15:0] a;
    reg [15:0] b;
    wire [15:0] out;

    Or16 mymodule(out, a, b);
    
    initial
    begin
        $dumpfile("tb_Or16.vcd");
        $dumpvars(0, tb_Or16);

        a = 16'b0000010001101010; b = 16'b1101111001010111; #1;
         `assert(out, 16'b1101111001111111)
        a = 16'b0000011111011000; b = 16'b0001000110011000; #1;
         `assert(out, 16'b0001011111011000)
        a = 16'b0001000011000000; b = 16'b1101011101101011; #1;
         `assert(out, 16'b1101011111101011)
        a = 16'b0001011010000101; b = 16'b0000110101000001; #1;
         `assert(out, 16'b0001111111000101)
        a = 16'b0001110111001011; b = 16'b1101101001100110; #1;
         `assert(out, 16'b1101111111101111)
        a = 16'b0010001011010110; b = 16'b0000101101001011; #1;
         `assert(out, 16'b0010101111011111)
        a = 16'b0010010101100010; b = 16'b0011100101011100; #1;
         `assert(out, 16'b0011110101111110)
        a = 16'b0010110100111001; b = 16'b1001100001111001; #1;
         `assert(out, 16'b1011110101111001)
        a = 16'b0010111100101110; b = 16'b1111011011011000; #1;
         `assert(out, 16'b1111111111111110)
        a = 16'b0011000100101110; b = 16'b0101001011101100; #1;
         `assert(out, 16'b0111001111101110)
        a = 16'b0011001010111100; b = 16'b0010001101100111; #1;
         `assert(out, 16'b0011001111111111)
        a = 16'b0011001101110010; b = 16'b1110000110100110; #1;
         `assert(out, 16'b1111001111110110)
        a = 16'b0100101100010001; b = 16'b1111111010001110; #1;
         `assert(out, 16'b1111111110011111)
        a = 16'b0101001000011011; b = 16'b0010001011011011; #1;
         `assert(out, 16'b0111001011011011)
        a = 16'b0101001101010100; b = 16'b1000100001010010; #1;
         `assert(out, 16'b1101101101010110)
        a = 16'b0101011101101011; b = 16'b0100000100110111; #1;
         `assert(out, 16'b0101011101111111)
        a = 16'b0111010100111111; b = 16'b1000010010100101; #1;
         `assert(out, 16'b1111010110111111)
        a = 16'b0111101111110110; b = 16'b1011111101010000; #1;
         `assert(out, 16'b1111111111110110)
        a = 16'b0111110111101111; b = 16'b1010110000001110; #1;
         `assert(out, 16'b1111110111101111)
        a = 16'b1000011111011101; b = 16'b0001111101101011; #1;
         `assert(out, 16'b1001111111111111)
        a = 16'b1000110000010011; b = 16'b0100101111100001; #1;
         `assert(out, 16'b1100111111110011)
        a = 16'b1000110101011001; b = 16'b0011001000010011; #1;
         `assert(out, 16'b1011111101011011)
        a = 16'b1001011001001000; b = 16'b0111110101101110; #1;
         `assert(out, 16'b1111111101101110)
        a = 16'b1001101011110111; b = 16'b1000100111101100; #1;
         `assert(out, 16'b1001101111111111)
        a = 16'b1010101000000010; b = 16'b0111001011000110; #1;
         `assert(out, 16'b1111101011000110)
        a = 16'b1011001100111001; b = 16'b0111001001011111; #1;
         `assert(out, 16'b1111001101111111)
        a = 16'b1011101011000001; b = 16'b1110001000010101; #1;
         `assert(out, 16'b1111101011010101)
        a = 16'b1100110111011000; b = 16'b0001000101101000; #1;
         `assert(out, 16'b1101110111111000)
        a = 16'b1100111001100101; b = 16'b1010010100110110; #1;
         `assert(out, 16'b1110111101110111)
        a = 16'b1111000111011001; b = 16'b1011000111000101; #1;
         `assert(out, 16'b1111000111011101)

    end
endmodule