/* testbench para RAM32 */
/* ordem de portas: out, in, addr, write, clk */
/* input [15:0] in; */
/* input [4:0] addr; */
/* input write, clk; */
/* output [15:0] out; */

`include "RAM32.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_RAM32;
    reg [15:0] in;
    reg [4:0] addr;
    reg write, clk;
    wire [15:0] out;

    RAM32 ram0(out, in, addr, write, clk);
    
    always
    begin
        #1 clk = ~clk;
    end
    
    initial
    begin
        $dumpfile("tb_RAM32.vcd");
        $dumpvars(0, tb_RAM32);

        clk = 0;

        /* Inicializa a memória zerando todos os registradores */
        in = 16'b0000000000000000; addr = 5'b00000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b00111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b01111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b10111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11111; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11000; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11001; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11010; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11011; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11100; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11101; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11110; write = 1; #3;
        in = 16'b0000000000000000; addr = 5'b11111; write = 1; #3;

        /* Testando leitura e escrita */
        in = 16'b0000000001110000; addr = 5'b00000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 5'b00001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 5'b00010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 5'b00011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 5'b00100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 5'b00101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 5'b00110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 5'b00111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 5'b00000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 5'b00001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 5'b00010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 5'b00011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 5'b00100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 5'b00101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 5'b00110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 5'b00111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 5'b00000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 5'b00001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 5'b00010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 5'b00011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 5'b00100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 5'b00101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 5'b00110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 5'b00111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 5'b01000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 5'b01001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 5'b01010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 5'b01011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 5'b01100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 5'b01101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 5'b01110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 5'b01111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 5'b01000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 5'b01001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 5'b01010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 5'b01011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 5'b01100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 5'b01101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 5'b01110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 5'b01111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 5'b01000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 5'b01001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 5'b01010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 5'b01011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 5'b01100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 5'b01101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 5'b01110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 5'b01111; write = 0; #3;
        `assert(out, 16'b0000000001110010);
    
        in = 16'b0000000001110000; addr = 5'b10000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 5'b10001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 5'b10010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 5'b10011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 5'b10100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 5'b10101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 5'b10110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 5'b10111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 5'b10000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 5'b10001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 5'b10010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 5'b10011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 5'b10100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 5'b10101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 5'b10110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 5'b10111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 5'b10000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 5'b10001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 5'b10010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 5'b10011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 5'b10100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 5'b10101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 5'b10110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 5'b10111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 5'b11000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 5'b11001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 5'b11010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 5'b11011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 5'b11100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 5'b11101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 5'b11110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 5'b11111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 5'b11000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 5'b11001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 5'b11010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 5'b11011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 5'b11100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 5'b11101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 5'b11110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 5'b11111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 5'b11000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 5'b11001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 5'b11010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 5'b11011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 5'b11100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 5'b11101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 5'b11110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 5'b11111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        $finish;
    end

endmodule
