/* testbench para DMux16 */
/* ordem de portas: a, b, in, sel */
/* input [15:0] in; input sel; */
/* output [15:0] a; output [15:0] b; */

`include "DMux16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_DMux16;
    reg [15:0] in;
    reg sel;
    wire [15:0] a;
    wire [15:0] b;

    DMux16 mymodule(a, b, in, sel);
    
    initial
    begin
        $dumpfile("tb_DMux16.vcd");
        $dumpvars(0, tb_DMux16);

        in = 16'b0000100100011110; sel = 1'b0; #1;
         `assert(a, 16'b0000100100011110) `assert(b, 16'b0000000000000000)
        in = 16'b0000110101100101; sel = 1'b0; #1;
         `assert(a, 16'b0000110101100101) `assert(b, 16'b0000000000000000)
        in = 16'b0001010110000000; sel = 1'b0; #1;
         `assert(a, 16'b0001010110000000) `assert(b, 16'b0000000000000000)
        in = 16'b0001010110111110; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0001010110111110)
        in = 16'b0001100010000011; sel = 1'b0; #1;
         `assert(a, 16'b0001100010000011) `assert(b, 16'b0000000000000000)
        in = 16'b0010000011110001; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0010000011110001)
        in = 16'b0010000100111011; sel = 1'b0; #1;
         `assert(a, 16'b0010000100111011) `assert(b, 16'b0000000000000000)
        in = 16'b0010010001110000; sel = 1'b0; #1;
         `assert(a, 16'b0010010001110000) `assert(b, 16'b0000000000000000)
        in = 16'b0010111110101011; sel = 1'b0; #1;
         `assert(a, 16'b0010111110101011) `assert(b, 16'b0000000000000000)
        in = 16'b0011111011000000; sel = 1'b0; #1;
         `assert(a, 16'b0011111011000000) `assert(b, 16'b0000000000000000)
        in = 16'b0100000000011100; sel = 1'b0; #1;
         `assert(a, 16'b0100000000011100) `assert(b, 16'b0000000000000000)
        in = 16'b0100100111011000; sel = 1'b0; #1;
         `assert(a, 16'b0100100111011000) `assert(b, 16'b0000000000000000)
        in = 16'b0101001110011111; sel = 1'b0; #1;
         `assert(a, 16'b0101001110011111) `assert(b, 16'b0000000000000000)
        in = 16'b0101011010110110; sel = 1'b0; #1;
         `assert(a, 16'b0101011010110110) `assert(b, 16'b0000000000000000)
        in = 16'b0101100110011000; sel = 1'b0; #1;
         `assert(a, 16'b0101100110011000) `assert(b, 16'b0000000000000000)
        in = 16'b0110101001010100; sel = 1'b0; #1;
         `assert(a, 16'b0110101001010100) `assert(b, 16'b0000000000000000)
        in = 16'b0110110100001000; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0110110100001000)
        in = 16'b1001001000111100; sel = 1'b0; #1;
         `assert(a, 16'b1001001000111100) `assert(b, 16'b0000000000000000)
        in = 16'b1001011101000101; sel = 1'b0; #1;
         `assert(a, 16'b1001011101000101) `assert(b, 16'b0000000000000000)
        in = 16'b1001111111001100; sel = 1'b0; #1;
         `assert(a, 16'b1001111111001100) `assert(b, 16'b0000000000000000)
        in = 16'b1010010011101000; sel = 1'b0; #1;
         `assert(a, 16'b1010010011101000) `assert(b, 16'b0000000000000000)
        in = 16'b1010011010100111; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1010011010100111)
        in = 16'b1100110001011111; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1100110001011111)
        in = 16'b1101011101100011; sel = 1'b0; #1;
         `assert(a, 16'b1101011101100011) `assert(b, 16'b0000000000000000)
        in = 16'b1101100010010000; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1101100010010000)
        in = 16'b1101111010001011; sel = 1'b0; #1;
         `assert(a, 16'b1101111010001011) `assert(b, 16'b0000000000000000)
        in = 16'b1110011001000110; sel = 1'b0; #1;
         `assert(a, 16'b1110011001000110) `assert(b, 16'b0000000000000000)
        in = 16'b1110100110111011; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1110100110111011)
        in = 16'b1111000000010000; sel = 1'b0; #1;
         `assert(a, 16'b1111000000010000) `assert(b, 16'b0000000000000000)
        in = 16'b1111000100100000; sel = 1'b1; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1111000100100000)

    end
endmodule