/* testbench para Mux8Way16 */
/* ordem de portas: out, a, b, c, d, e, f, g, h, sel */
/* input [15:0] a; input [15:0] b; input [15:0] c; input [15:0] d; input [15:0] e; input [15:0] f; input [15:0] g; input [15:0] h; input [2:0] sel; */
/* output [15:0] out; */

`include "Mux8Way16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_Mux8Way16;
    reg [15:0] a;
    reg [15:0] b;
    reg [15:0] c;
    reg [15:0] d;
    reg [15:0] e;
    reg [15:0] f;
    reg [15:0] g;
    reg [15:0] h;
    reg [2:0] sel;
    wire [15:0] out;

    Mux8Way16 mymodule(out, a, b, c, d, e, f, g, h, sel);
    
    initial
    begin
        $dumpfile("tb_Mux8Way16.vcd");
        $dumpvars(0, tb_Mux8Way16);

        a = 16'b0000000000000000; b = 16'b0000000000000000; c = 16'b0000000000000000; d = 16'b0000000000000000; e = 16'b0000000000000000; f = 16'b0000000000000000; g = 16'b0000000000000000; h = 16'b0000000000000000; sel = 3'b000; #1;
         `assert(out, 16'b0000000000000000)
        a = 16'b0001001000100111; b = 16'b0110100001010001; c = 16'b0011110000010100; d = 16'b1111111111011000; e = 16'b1100010000110101; f = 16'b0111101000101001; g = 16'b1001010101100000; h = 16'b1101101000101100; sel = 3'b111; #1;
         `assert(out, 16'b1101101000101100)
        a = 16'b0001100100111000; b = 16'b0101011100111110; c = 16'b1101011000101010; d = 16'b0000001101011100; e = 16'b0010101100101000; f = 16'b1110011010110011; g = 16'b0111111001000110; h = 16'b0000110010010100; sel = 3'b000; #1;
         `assert(out, 16'b0001100100111000)
        a = 16'b0010110110111011; b = 16'b1010101001000000; c = 16'b1010011011101100; d = 16'b0000100011100011; e = 16'b1101110110011111; f = 16'b1100111001000111; g = 16'b1010010000011000; h = 16'b1110001101010101; sel = 3'b110; #1;
         `assert(out, 16'b1010010000011000)
        a = 16'b0011000011011001; b = 16'b0011110001101010; c = 16'b1110011111011000; d = 16'b0000100010110100; e = 16'b1110101010011000; f = 16'b0001010100101110; g = 16'b1100111110110000; h = 16'b1010011100100010; sel = 3'b111; #1;
         `assert(out, 16'b1010011100100010)
        a = 16'b0011101011111010; b = 16'b0010010011111100; c = 16'b0010100101100110; d = 16'b1001000100100010; e = 16'b0000010001011010; f = 16'b0001010011011100; g = 16'b0001111110100001; h = 16'b1111001011011001; sel = 3'b100; #1;
         `assert(out, 16'b0000010001011010)
        a = 16'b0100011001010100; b = 16'b1010101001010111; c = 16'b1111011110010110; d = 16'b1000101100010110; e = 16'b1110110010000101; f = 16'b1001100000111000; g = 16'b1111101100110110; h = 16'b1001111000011010; sel = 3'b001; #1;
         `assert(out, 16'b1010101001010111)
        a = 16'b0100110000000111; b = 16'b1111001111100111; c = 16'b1001000100111010; d = 16'b0000001011111110; e = 16'b1110011010000110; f = 16'b0001101110111001; g = 16'b0111111111101011; h = 16'b1110111001110100; sel = 3'b010; #1;
         `assert(out, 16'b1001000100111010)
        a = 16'b0100111110011100; b = 16'b0011110101000011; c = 16'b1100101111101110; d = 16'b0011010011001010; e = 16'b1100110001001010; f = 16'b0010000011000101; g = 16'b1010100001111010; h = 16'b0010011100000010; sel = 3'b000; #1;
         `assert(out, 16'b0100111110011100)
        a = 16'b0101000010111111; b = 16'b0000001011110000; c = 16'b0110100010101011; d = 16'b0101101001000100; e = 16'b1100000001101001; f = 16'b0011011111100101; g = 16'b0001010010000111; h = 16'b1111001111100100; sel = 3'b000; #1;
         `assert(out, 16'b0101000010111111)
        a = 16'b0110001101110001; b = 16'b0010111110000100; c = 16'b0111111110110101; d = 16'b1010100001100100; e = 16'b1110010111001101; f = 16'b1110100111101100; g = 16'b1111000101011010; h = 16'b0100011110111101; sel = 3'b011; #1;
         `assert(out, 16'b1010100001100100)
        a = 16'b0110111010110100; b = 16'b1111010110101100; c = 16'b0101000001110111; d = 16'b1011010001101100; e = 16'b1011110010110010; f = 16'b0110010100010011; g = 16'b0000111100111011; h = 16'b1001100110101010; sel = 3'b000; #1;
         `assert(out, 16'b0110111010110100)
        a = 16'b0111001111010101; b = 16'b0011011000110000; c = 16'b1111111000011100; d = 16'b1000011001000101; e = 16'b1010010101000110; f = 16'b0011101010010011; g = 16'b1001010000110000; h = 16'b0010011110100011; sel = 3'b001; #1;
         `assert(out, 16'b0011011000110000)
        a = 16'b1000001111110001; b = 16'b1101100101011111; c = 16'b1011100001101101; d = 16'b0001100010010100; e = 16'b1001111001011011; f = 16'b1101001011010010; g = 16'b1000010000111001; h = 16'b1011110001101010; sel = 3'b000; #1;
         `assert(out, 16'b1000001111110001)
        a = 16'b1000010111110001; b = 16'b1110110110100000; c = 16'b1011010010010001; d = 16'b1011000100010110; e = 16'b1001100011001010; f = 16'b0001100101010110; g = 16'b0101010001111110; h = 16'b1000100111101101; sel = 3'b100; #1;
         `assert(out, 16'b1001100011001010)
        a = 16'b1010010000011110; b = 16'b0011101000010011; c = 16'b1010010011001000; d = 16'b0100111000100111; e = 16'b0101001100101001; f = 16'b0100001000111000; g = 16'b1001101001111101; h = 16'b0011100010100011; sel = 3'b010; #1;
         `assert(out, 16'b1010010011001000)
        a = 16'b1010011011101101; b = 16'b1101101011101111; c = 16'b0000101010011001; d = 16'b1111001011011100; e = 16'b1010010000000100; f = 16'b1101101110000010; g = 16'b1010010110011101; h = 16'b1010110000011111; sel = 3'b000; #1;
         `assert(out, 16'b1010011011101101)
        a = 16'b1011001101000101; b = 16'b0000010000010111; c = 16'b0011101010000000; d = 16'b0010000010101111; e = 16'b1001101010111000; f = 16'b0001001011011110; g = 16'b1110100001010100; h = 16'b0001111010001000; sel = 3'b101; #1;
         `assert(out, 16'b0001001011011110)
        a = 16'b1011100111100010; b = 16'b0100000111100110; c = 16'b0111000000100100; d = 16'b0101000110001101; e = 16'b0011111011110111; f = 16'b1000101000111000; g = 16'b0111110001001001; h = 16'b1111001110111101; sel = 3'b000; #1;
         `assert(out, 16'b1011100111100010)
        a = 16'b1011111101100000; b = 16'b0010010100011111; c = 16'b0110000010101111; d = 16'b0001001010010110; e = 16'b0010010011000110; f = 16'b0011001000010010; g = 16'b1101111111101101; h = 16'b1000111111100000; sel = 3'b001; #1;
         `assert(out, 16'b0010010100011111)
        a = 16'b1100000010000111; b = 16'b1000000111000011; c = 16'b0101111111000010; d = 16'b0100000010101011; e = 16'b0010101011010010; f = 16'b0101100100010000; g = 16'b0011110010101100; h = 16'b1011111010101110; sel = 3'b000; #1;
         `assert(out, 16'b1100000010000111)
        a = 16'b1100010100010011; b = 16'b0101111010111010; c = 16'b0000010111101110; d = 16'b0000110100110001; e = 16'b1010101000111100; f = 16'b0011011111110100; g = 16'b0011011100000111; h = 16'b1100111100101001; sel = 3'b100; #1;
         `assert(out, 16'b1010101000111100)
        a = 16'b1100011110111010; b = 16'b1110101110110001; c = 16'b1000011100110111; d = 16'b1001111010010110; e = 16'b1101011101011000; f = 16'b0101011110110101; g = 16'b0010100101000011; h = 16'b0010011101001100; sel = 3'b110; #1;
         `assert(out, 16'b0010100101000011)
        a = 16'b1101000001100111; b = 16'b1111111000011011; c = 16'b1011000010110000; d = 16'b0100111000101001; e = 16'b0100100010100010; f = 16'b0110100110000111; g = 16'b1000011000011100; h = 16'b1010111110010111; sel = 3'b101; #1;
         `assert(out, 16'b0110100110000111)
        a = 16'b1101101001000000; b = 16'b1100010001111011; c = 16'b0110111110011101; d = 16'b0111101001110011; e = 16'b1110011110010110; f = 16'b0111111000010100; g = 16'b1100010010010011; h = 16'b0111010101110001; sel = 3'b011; #1;
         `assert(out, 16'b0111101001110011)
        a = 16'b1110110111110101; b = 16'b1001011111011000; c = 16'b1101010111011100; d = 16'b0100000100010001; e = 16'b0111110001010000; f = 16'b0110110101101011; g = 16'b0110010111101100; h = 16'b1110011011111101; sel = 3'b111; #1;
         `assert(out, 16'b1110011011111101)
        a = 16'b1110111110000101; b = 16'b0111101000111111; c = 16'b1011001100100111; d = 16'b1111000011101100; e = 16'b0101001011100000; f = 16'b1111101011111001; g = 16'b0010001011001110; h = 16'b1000110000011011; sel = 3'b110; #1;
         `assert(out, 16'b0010001011001110)
        a = 16'b1111101001010101; b = 16'b1010001101100011; c = 16'b0000000100000101; d = 16'b0101100011101011; e = 16'b0001101111100010; f = 16'b0100101011000110; g = 16'b1011011101001001; h = 16'b1011011111010110; sel = 3'b010; #1;
         `assert(out, 16'b0000000100000101)
        a = 16'b1111110100000100; b = 16'b1011000101100010; c = 16'b0010000101111010; d = 16'b1110011110100100; e = 16'b0010010011001010; f = 16'b0001000001010001; g = 16'b0000101101101100; h = 16'b0011000000001101; sel = 3'b011; #1;
         `assert(out, 16'b1110011110100100)
        a = 16'b1111111111111111; b = 16'b1111111111111111; c = 16'b1111111111111111; d = 16'b1111111111111111; e = 16'b1111111111111111; f = 16'b1111111111111111; g = 16'b1111111111111111; h = 16'b1111111111111111; sel = 3'b111; #1;
         `assert(out, 16'b1111111111111111)

    end
endmodule