/* testbench para DMux4Way16 */
/* ordem de portas: a, b, c, d, in, sel */
/* input [15:0] in; input [1:0] sel; */
/* output [15:0] a; output [15:0] b; output [15:0] c; output [15:0] d; */

`include "DMux4Way16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_DMux4Way16;
    reg [15:0] in;
    reg [1:0] sel;
    wire [15:0] a;
    wire [15:0] b;
    wire [15:0] c;
    wire [15:0] d;

    DMux4Way16 mymodule(a, b, c, d, in, sel);
    
    initial
    begin
        $dumpfile("tb_DMux4Way16.vcd");
        $dumpvars(0, tb_DMux4Way16);

        in = 16'b0000000000000000; sel = 2'b00; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0000001100111010; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000001100111010) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0000010000100110; sel = 2'b10; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000010000100110) `assert(d, 16'b0000000000000000)
        in = 16'b0001110110010111; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0001110110010111) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0010001101011001; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0010001101011001) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0010011111100000; sel = 2'b00; #1;
         `assert(a, 16'b0010011111100000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0010111000000001; sel = 2'b10; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0010111000000001) `assert(d, 16'b0000000000000000)
        in = 16'b0011100101100101; sel = 2'b10; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0011100101100101) `assert(d, 16'b0000000000000000)
        in = 16'b0011110011001111; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0011110011001111)
        in = 16'b0100100110100000; sel = 2'b00; #1;
         `assert(a, 16'b0100100110100000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0100111010101010; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0100111010101010) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0101100000100110; sel = 2'b00; #1;
         `assert(a, 16'b0101100000100110) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0101111110101101; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0101111110101101)
        in = 16'b0110101110110101; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0110101110110101) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b0110111010011011; sel = 2'b10; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0110111010011011) `assert(d, 16'b0000000000000000)
        in = 16'b0111111100110111; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0111111100110111)
        in = 16'b1000000110001110; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1000000110001110)
        in = 16'b1000001110110011; sel = 2'b10; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b1000001110110011) `assert(d, 16'b0000000000000000)
        in = 16'b1001010100111000; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1001010100111000)
        in = 16'b1010011010110100; sel = 2'b00; #1;
         `assert(a, 16'b1010011010110100) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b1010111111001101; sel = 2'b00; #1;
         `assert(a, 16'b1010111111001101) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b1011101000110011; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1011101000110011)
        in = 16'b1100000000101001; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1100000000101001) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b1101001111110111; sel = 2'b00; #1;
         `assert(a, 16'b1101001111110111) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b1101010000110001; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1101010000110001) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b1110000010001010; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1110000010001010)
        in = 16'b1110001110010101; sel = 2'b01; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b1110001110010101) `assert(c, 16'b0000000000000000) `assert(d, 16'b0000000000000000)
        in = 16'b1111011111000000; sel = 2'b10; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b1111011111000000) `assert(d, 16'b0000000000000000)
        in = 16'b1111110010110001; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1111110010110001)
        in = 16'b1111111111111111; sel = 2'b11; #1;
         `assert(a, 16'b0000000000000000) `assert(b, 16'b0000000000000000) `assert(c, 16'b0000000000000000) `assert(d, 16'b1111111111111111)

    end
endmodule