/* testbench para And16 */
/* ordem de portas: out, a, b */
/* input [15:0] a; input [15:0] b; */
/* output [15:0] out; */

`include "And16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_And16;
    reg [15:0] a;
    reg [15:0] b;
    wire [15:0] out;

    And16 mymodule(out, a, b);
    
    initial
    begin
        $dumpfile("tb_And16.vcd");
        $dumpvars(0, tb_And16);

        a = 16'b0000001101110001; b = 16'b1100111011100000; #1;
         `assert(out, 16'b0000001001100000)
        a = 16'b0000010000101011; b = 16'b0110110100101110; #1;
         `assert(out, 16'b0000010000101010)
        a = 16'b0000101000110001; b = 16'b1010001001110001; #1;
         `assert(out, 16'b0000001000110001)
        a = 16'b0000101100110110; b = 16'b1011101001110101; #1;
         `assert(out, 16'b0000101000110100)
        a = 16'b0001010000011111; b = 16'b1111101101011001; #1;
         `assert(out, 16'b0001000000011001)
        a = 16'b0001010000100010; b = 16'b1010000110001100; #1;
         `assert(out, 16'b0000000000000000)
        a = 16'b0001101001101000; b = 16'b1010001011100110; #1;
         `assert(out, 16'b0000001001100000)
        a = 16'b0001110111010011; b = 16'b0000101010101100; #1;
         `assert(out, 16'b0000100010000000)
        a = 16'b0010011000100110; b = 16'b1001001000100101; #1;
         `assert(out, 16'b0000001000100100)
        a = 16'b0010111011101000; b = 16'b0111101001111100; #1;
         `assert(out, 16'b0010101001101000)
        a = 16'b0100010110001111; b = 16'b0100011010111110; #1;
         `assert(out, 16'b0100010010001110)
        a = 16'b0100010110100011; b = 16'b1001110100111100; #1;
         `assert(out, 16'b0000010100100000)
        a = 16'b0100110010011111; b = 16'b0111011111100000; #1;
         `assert(out, 16'b0100010010000000)
        a = 16'b0100111011000011; b = 16'b0100101100000011; #1;
         `assert(out, 16'b0100101000000011)
        a = 16'b0101111001100000; b = 16'b0100000010011001; #1;
         `assert(out, 16'b0100000000000000)
        a = 16'b0110000001111010; b = 16'b0000100001011111; #1;
         `assert(out, 16'b0000000001011010)
        a = 16'b0110000011110011; b = 16'b1100001000001111; #1;
         `assert(out, 16'b0100000000000011)
        a = 16'b0110010101001101; b = 16'b0110100001011101; #1;
         `assert(out, 16'b0110000001001101)
        a = 16'b0111000101110001; b = 16'b0111001001000110; #1;
         `assert(out, 16'b0111000001000000)
        a = 16'b0111100110011100; b = 16'b0101110010100011; #1;
         `assert(out, 16'b0101100010000000)
        a = 16'b1000010110010100; b = 16'b0000000111010001; #1;
         `assert(out, 16'b0000000110010000)
        a = 16'b1001001100101110; b = 16'b0100100000100010; #1;
         `assert(out, 16'b0000000000100010)
        a = 16'b1001101111101110; b = 16'b1000011111110001; #1;
         `assert(out, 16'b1000001111100000)
        a = 16'b1010100110010000; b = 16'b1000111011000100; #1;
         `assert(out, 16'b1000100010000000)
        a = 16'b1011110010100100; b = 16'b0100000010100111; #1;
         `assert(out, 16'b0000000010100100)
        a = 16'b1100100000010001; b = 16'b1001110100111110; #1;
         `assert(out, 16'b1000100000010000)
        a = 16'b1100100101111010; b = 16'b1011001110000001; #1;
         `assert(out, 16'b1000000100000000)
        a = 16'b1101001100011000; b = 16'b1111011010100100; #1;
         `assert(out, 16'b1101001000000000)
        a = 16'b1110101110100000; b = 16'b1111011100101101; #1;
         `assert(out, 16'b1110001100100000)
        a = 16'b1111111111111101; b = 16'b0100110100101101; #1;
         `assert(out, 16'b0100110100101101)

    end
endmodule