/* testbench para Mux4Way16 */
/* ordem de portas: out, a, b, c, d, sel */
/* input [15:0] a; input [15:0] b; input [15:0] c; input [15:0] d; input [1:0] sel; */
/* output [15:0] out; */

`include "Mux4Way16.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_Mux4Way16;
    reg [15:0] a;
    reg [15:0] b;
    reg [15:0] c;
    reg [15:0] d;
    reg [1:0] sel;
    wire [15:0] out;

    Mux4Way16 mymodule(out, a, b, c, d, sel);
    
    initial
    begin
        $dumpfile("tb_Mux4Way16.vcd");
        $dumpvars(0, tb_Mux4Way16);

        a = 16'b0000000000000000; b = 16'b0000000000000000; c = 16'b0000000000000000; d = 16'b0000000000000000; sel = 2'b00; #1;
         `assert(out, 16'b0000000000000000)
        a = 16'b1110000111011000; b = 16'b0110001001111011; c = 16'b0110000101001011; d = 16'b1001110010010011; sel = 2'b01; #1;
         `assert(out, 16'b0110001001111011)
        a = 16'b1110100010010010; b = 16'b0101111000001000; c = 16'b1100010110110111; d = 16'b0011011010100011; sel = 2'b01; #1;
         `assert(out, 16'b0101111000001000)
        a = 16'b1110100101111000; b = 16'b1100011100111001; c = 16'b0000011100010010; d = 16'b1101100011111101; sel = 2'b00; #1;
         `assert(out, 16'b1110100101111000)
        a = 16'b1110101011000101; b = 16'b0110110001101000; c = 16'b1000011011100000; d = 16'b1101001111010100; sel = 2'b01; #1;
         `assert(out, 16'b0110110001101000)
        a = 16'b1110110001100011; b = 16'b1010111111000111; c = 16'b1100111000100001; d = 16'b1110011001001000; sel = 2'b10; #1;
         `assert(out, 16'b1100111000100001)
        a = 16'b1111000101111100; b = 16'b1000011101101010; c = 16'b0110001110000001; d = 16'b1001101001010101; sel = 2'b00; #1;
         `assert(out, 16'b1111000101111100)
        a = 16'b1111001010011110; b = 16'b1100000100011101; c = 16'b1011101110110101; d = 16'b0110101111011110; sel = 2'b10; #1;
         `assert(out, 16'b1011101110110101)
        a = 16'b1111001011000101; b = 16'b0100101000010000; c = 16'b1001011110011110; d = 16'b1101111110001111; sel = 2'b10; #1;
         `assert(out, 16'b1001011110011110)
        a = 16'b1111001100110100; b = 16'b0011110100110000; c = 16'b0110001100111011; d = 16'b0101100000010010; sel = 2'b11; #1;
         `assert(out, 16'b0101100000010010)
        a = 16'b1111001110001000; b = 16'b1101011000100011; c = 16'b1101011011110101; d = 16'b1001000111001001; sel = 2'b11; #1;
         `assert(out, 16'b1001000111001001)
        a = 16'b1111100110011011; b = 16'b0110111111001110; c = 16'b1001001000011000; d = 16'b1000110010000101; sel = 2'b01; #1;
         `assert(out, 16'b0110111111001110)
        a = 16'b1111101101001100; b = 16'b1001100111011010; c = 16'b0010011000110110; d = 16'b1111110101001110; sel = 2'b01; #1;
         `assert(out, 16'b1001100111011010)
        a = 16'b1111111001111111; b = 16'b0111100110001000; c = 16'b0111110100011000; d = 16'b0000101000110000; sel = 2'b11; #1;
         `assert(out, 16'b0000101000110000)
        a = 16'b0000001000111101; b = 16'b1110011111001100; c = 16'b1110010111001110; d = 16'b0001001001011101; sel = 2'b10; #1;
         `assert(out, 16'b1110010111001110)
        a = 16'b0000001011110011; b = 16'b1101101010100001; c = 16'b0110111100101010; d = 16'b0100110001000110; sel = 2'b01; #1;
         `assert(out, 16'b1101101010100001)
        a = 16'b0000010001011100; b = 16'b0110000101000111; c = 16'b0010100111100100; d = 16'b1111001010011100; sel = 2'b11; #1;
         `assert(out, 16'b1111001010011100)
        a = 16'b0000011001010000; b = 16'b0011000110010011; c = 16'b0111010110000010; d = 16'b0011010111011010; sel = 2'b11; #1;
         `assert(out, 16'b0011010111011010)
        a = 16'b0000011110100110; b = 16'b0100110111011011; c = 16'b0000101100000100; d = 16'b0101010100111000; sel = 2'b01; #1;
         `assert(out, 16'b0100110111011011)
        a = 16'b0000100011101101; b = 16'b0111100001111100; c = 16'b0011110011011010; d = 16'b0110011000010001; sel = 2'b01; #1;
         `assert(out, 16'b0111100001111100)
        a = 16'b0000101011001111; b = 16'b1110110110100001; c = 16'b1010001111000010; d = 16'b0111001000010100; sel = 2'b11; #1;
         `assert(out, 16'b0111001000010100)
        a = 16'b0000110001001110; b = 16'b1111100101001011; c = 16'b0010011100011111; d = 16'b0100110010010101; sel = 2'b10; #1;
         `assert(out, 16'b0010011100011111)
        a = 16'b0000110010110001; b = 16'b1110000011001001; c = 16'b1011010100100011; d = 16'b1111100111100110; sel = 2'b10; #1;
         `assert(out, 16'b1011010100100011)
        a = 16'b0001010011010001; b = 16'b0011001110111010; c = 16'b0010111001000011; d = 16'b1010001100100010; sel = 2'b10; #1;
         `assert(out, 16'b0010111001000011)
        a = 16'b0001011010001001; b = 16'b1000000111000100; c = 16'b0100011011001010; d = 16'b1010100000100110; sel = 2'b01; #1;
         `assert(out, 16'b1000000111000100)
        a = 16'b0001011101110111; b = 16'b1010101010011101; c = 16'b1100110101000100; d = 16'b1001100010100001; sel = 2'b01; #1;
         `assert(out, 16'b1010101010011101)
        a = 16'b0001111000010110; b = 16'b0001000010111111; c = 16'b1110010010000110; d = 16'b1100001111011110; sel = 2'b10; #1;
         `assert(out, 16'b1110010010000110)
        a = 16'b0001111001000011; b = 16'b0110110111000001; c = 16'b1101000011011100; d = 16'b1111010101111100; sel = 2'b00; #1;
         `assert(out, 16'b0001111001000011)
        a = 16'b0001111010011011; b = 16'b0100011010000000; c = 16'b1111101101010000; d = 16'b0110111111000101; sel = 2'b11; #1;
         `assert(out, 16'b0110111111000101)
        a = 16'b1111111111111111; b = 16'b1111111111111111; c = 16'b1111111111111111; d = 16'b1111111111111111; sel = 2'b11; #1;
         `assert(out, 16'b1111111111111111)

    end
endmodule