/* testbench para RAM64 */
/* ordem de portas: out, in, addr, write, clk */
/* input [15:0] in; */
/* input [4:0] addr; */
/* input write, clk; */
/* output [15:0] out; */

`include "RAM64.v"

`define assert(signal, value) \
    if (signal !== value) \
    begin \
        $display("ASSERTION FAILED in %m: signal != value"); \
        $finish; \
    end else begin \
        $display("Success! %m: signal = value"); \
    end

module tb_RAM64;
    reg [15:0] in;
    reg [5:0] addr;
    reg write, clk;
    wire [15:0] out;

    RAM64 ram0(out, in, addr, write, clk);
    
    always
    begin
        #1 clk = ~clk;
    end
    
    initial
    begin
        $dumpfile("tb_RAM64.vcd");
        $dumpvars(0, tb_RAM64);

        clk = 0;

        /* Inicializa a memória zerando todos os registradores */
        in = 16'b0000000000000000; addr = 6'b000000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b000111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b001111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b010111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b011111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b100111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b101111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b110111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111111; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111000; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111001; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111010; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111011; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111100; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111101; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111110; write = 1; #3;
        in = 16'b0000000000000000; addr = 6'b111111; write = 1; #3;

        /* Testando leitura e escrita */
        in = 16'b0000000001110000; addr = 6'b000000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b000001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b000010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b000011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b000100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b000101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b000110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b000111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b000000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b000001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b000010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b000011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b000100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b000101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b000110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b000111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b000000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b000001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b000010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b000011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b000100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b000101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b000110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b000111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 6'b001000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b001001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b001010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b001011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b001100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b001101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b001110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b001111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b001000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b001001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b001010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b001011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b001100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b001101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b001110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b001111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b001000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b001001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b001010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b001011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b001100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b001101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b001110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b001111; write = 0; #3;
        `assert(out, 16'b0000000001110010);
    
        in = 16'b0000000001110000; addr = 6'b010000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b010001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b010010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b010011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b010100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b010101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b010110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b010111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b010000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b010001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b010010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b010011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b010100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b010101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b010110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b010111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b010000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b010001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b010010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b010011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b010100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b010101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b010110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b010111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 6'b011000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b011001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b011010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b011011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b011100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b011101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b011110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b011111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b011000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b011001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b011010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b011011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b011100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b011101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b011110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b011111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b011000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b011001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b011010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b011011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b011100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b011101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b011110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b011111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 6'b100000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b100001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b100010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b100011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b100100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b100101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b100110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b100111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b100000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b100001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b100010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b100011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b100100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b100101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b100110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b100111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b100000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b100001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b100010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b100011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b100100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b100101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b100110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b100111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 6'b101000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b101001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b101010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b101011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b101100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b101101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b101110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b101111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b101000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b101001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b101010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b101011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b101100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b101101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b101110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b101111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b101000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b101001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b101010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b101011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b101100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b101101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b101110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b101111; write = 0; #3;
        `assert(out, 16'b0000000001110010);
    
        in = 16'b0000000001110000; addr = 6'b110000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b110001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b110010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b110011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b110100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b110101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b110110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b110111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b110000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b110001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b110010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b110011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b110100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b110101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b110110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b110111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b110000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b110001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b110010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b110011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b110100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b110101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b110110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b110111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000001110000; addr = 6'b111000; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100101; addr = 6'b111001; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100011; addr = 6'b111010; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110101; addr = 6'b111011; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101100; addr = 6'b111100; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001101001; addr = 6'b111101; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001100001; addr = 6'b111110; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110010; addr = 6'b111111; write = 0; #3;
        `assert(out, 16'b0000000000000000);

        in = 16'b0000000001110000; addr = 6'b111000; write = 1; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000001100101; addr = 6'b111001; write = 1; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000001100011; addr = 6'b111010; write = 1; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000001110101; addr = 6'b111011; write = 1; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000001101100; addr = 6'b111100; write = 1; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000001101001; addr = 6'b111101; write = 1; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000001100001; addr = 6'b111110; write = 1; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000001110010; addr = 6'b111111; write = 1; #3;
        `assert(out, 16'b0000000001110010);

        in = 16'b0000000000000000; addr = 6'b111000; write = 0; #3;
        `assert(out, 16'b0000000001110000);

        in = 16'b0000000000000000; addr = 6'b111001; write = 0; #3;
        `assert(out, 16'b0000000001100101);

        in = 16'b0000000000000000; addr = 6'b111010; write = 0; #3;
        `assert(out, 16'b0000000001100011);

        in = 16'b0000000000000000; addr = 6'b111011; write = 0; #3;
        `assert(out, 16'b0000000001110101);

        in = 16'b0000000000000000; addr = 6'b111100; write = 0; #3;
        `assert(out, 16'b0000000001101100);

        in = 16'b0000000000000000; addr = 6'b111101; write = 0; #3;
        `assert(out, 16'b0000000001101001);

        in = 16'b0000000000000000; addr = 6'b111110; write = 0; #3;
        `assert(out, 16'b0000000001100001);

        in = 16'b0000000000000000; addr = 6'b111111; write = 0; #3;
        `assert(out, 16'b0000000001110010);

        $finish;
    end

endmodule
